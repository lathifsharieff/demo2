module fifo (
    mod_name instance_name (.*);
    ports
);
    
endmodule